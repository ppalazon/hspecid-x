// `ifndef DATA_WIDTH
//   `define DATA_WIDTH 16
// `endif
// `ifndef DATA_WIDTH_MUL
//   `define DATA_WIDTH_MUL 32
// `endif
// `ifndef DATA_WIDTH_ACC
//   `define DATA_WIDTH_ACC 48
// `endif
// `ifndef VECTOR_LENGTH
//   `define VECTOR_LENGTH 24
// `endif
// `ifndef LENGTH_BITS
//   `define LENGTH_BITS 10
// `endif
// `ifndef BUFFER_LENGTH
//   `define BUFFER_LENGTH 4
// `endif
// `ifndef HSI_BANDS
//   `define HSI_BANDS 128
// `endif
