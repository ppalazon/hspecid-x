`timescale 1ns / 1ps

import hsid_pkg::*;
import ctrl_reg_tb_tasks::*;
import hsid_x_ctrl_reg_pkg::*;

module hsid_x_top_tb #(
    parameter WORD_WIDTH = HSID_WORD_WIDTH,  // Width of the word in bits
    parameter DATA_WIDTH_MUL = HSID_DATA_WIDTH_MUL,  // Data width for multiplication, larger than DATA_WIDTH
    parameter DATA_WIDTH_ACC = HSID_DATA_WIDTH_ACC,  // Data width for accumulator, larger than DATA_WIDTH
    parameter DATA_WIDTH = HSID_DATA_WIDTH,  // 16 bits by default
    parameter HSP_LIBRARY_WIDTH = HSID_HSP_LIBRARY_WIDTH,
    parameter HSP_BANDS_WIDTH = HSID_HSP_BANDS_WIDTH,
    parameter BUFFER_WIDTH = HSID_FIFO_ADDR_WIDTH,  // Length of the buffer
    parameter TEST_MEM_MASK = 32'h0000FFFF  // Mask to return least significant 14 bits of the address
  ) ();

  reg clk;
  reg rst_n;
  hsid_x_reg_pkg::reg_req_t reg_req;
  hsid_x_reg_pkg::reg_rsp_t reg_rsp;
  hsid_x_obi_inf_pkg::obi_resp_t obi_rsp;
  hsid_x_obi_inf_pkg::obi_req_t obi_req;
  wire hsid_x_int_o;

  reg random_gnt; // Random grant signal

  // Compute expected mse values for each pixel in the library
  logic [DATA_WIDTH-1:0] captured_hsp [];
  logic [DATA_WIDTH-1:0] reference_hsp [];
  logic [DATA_WIDTH_ACC:0] acc_int [];
  logic [WORD_WIDTH-1:0] expected_mse [];
  logic expected_mse_of [];
  logic [WORD_WIDTH-1:0] da_addr; // Direct access address
  logic [WORD_WIDTH-1:0] min_mse_value_expected;
  logic [WORD_WIDTH-1:0] max_mse_value_expected;
  logic [HSP_LIBRARY_WIDTH-1:0] min_mse_ref_expected;
  logic [HSP_LIBRARY_WIDTH-1:0] max_mse_ref_expected;

  hsid_x_top #(
    .WORD_WIDTH(WORD_WIDTH),
    .DATA_WIDTH(DATA_WIDTH),
    .DATA_WIDTH_MUL(DATA_WIDTH_MUL),
    .DATA_WIDTH_ACC(DATA_WIDTH_ACC),
    .BUFFER_WIDTH(BUFFER_WIDTH),
    .HSP_BANDS_WIDTH(HSP_BANDS_WIDTH),
    .HSP_LIBRARY_WIDTH(HSP_LIBRARY_WIDTH)
  ) dut (
    .clk(clk),
    .rst_n(rst_n),
    .reg_req_i(reg_req),
    .reg_rsp_o(reg_rsp),
    .obi_rsp_i(obi_rsp),
    .obi_req_o(obi_req),
    .hsid_x_int_o(hsid_x_int_o)
  );

  // Register interface debug
  reg_inf_debug reg_inf_debug_inst (
    .clk    (clk),
    .reg_req(reg_req),
    .reg_rsp(reg_rsp),
    .rst_n  (rst_n)
  );

  // OBI bus
  obi_bus_debug obi_bus_debug_inst (
    .clk    (clk),
    .rst_n  (rst_n),
    .obi_req(obi_req),
    .obi_rsp(obi_rsp)
  );

  // Connect test memory on the OBI bus
  pixel_obi_mem #(
    .DATA_WIDTH(DATA_WIDTH),
    .VALUE_MASK(TEST_MEM_MASK)
  ) u_pixel_obi_mem (
    .clk(clk),
    .rst_n(rst_n),
    .obi_req(obi_req),
    .obi_rsp(obi_rsp),
    .random_gnt(random_gnt)
  );

  const int STATUS_START = 32'b000001;
  const int STATUS_CLEAR = 32'b010000;
  const int STATUS_IDLE = 32'b000010;
  const int STATUS_DONE = 32'b001000;

  logic [WORD_WIDTH-1:0] library_size_w;
  logic [WORD_WIDTH-1:0] pixel_bands_w;
  logic [WORD_WIDTH-1:0] captured_pixel_addr_w;
  logic [WORD_WIDTH-1:0] library_pixel_addr_w;

  // Constrained randomization classes
  HsidXTopGen #(
    .WORD_WIDTH(WORD_WIDTH),
    .DATA_WIDTH(DATA_WIDTH),
    .DATA_WIDTH_MUL(DATA_WIDTH_MUL),  // Data width for multiplication, larger than DATA_WIDTH
    .DATA_WIDTH_ACC(DATA_WIDTH_ACC),  // Data width for accumulator, larger than DATA_WIDTH
    .HSP_BANDS_WIDTH(HSP_BANDS_WIDTH), // Address width for HSP bands
    .HSP_LIBRARY_WIDTH(HSP_LIBRARY_WIDTH) // Address width for HSI library
  ) hsid_x_top_gen = new();

  // Waveform generation for debugging
  initial begin
    $dumpfile("wave.vcd");
    $dumpvars(0, hsid_x_top_tb);
  end

  // Compute expected MSE values for each pixel in the library
  initial begin

    clk = 1;
    rst_n = 1;
    reg_req = hsid_x_reg_pkg::reg_req_t'(0);
    random_gnt = 0;

    #3 rst_n = 0; // Reset the DUT
    #5 rst_n = 1; // Release reset

    $display("Case 1: Normal scenario with constrained random cases...");
    for (int i = 0; i < 10; i++) begin
      if(!hsid_x_top_gen.randomize()) $fatal(0, "Randomization failed");

      // Get captured pixel data from the memory
      expected_pixel_mem(hsid_x_top_gen.captured_pixel_addr_w, hsid_x_top_gen.hsp_bands, captured_hsp);
      $display("Test %0d: Captured Pixel Address: 0x%0h, Library Address: 0x%0h, HSP Bands: %0d, Library size: %0d", i,
        hsid_x_top_gen.captured_pixel_addr_w, hsid_x_top_gen.library_pixel_addr_w, hsid_x_top_gen.hsp_bands, hsid_x_top_gen.library_size);
      hsid_x_top_gen.display_hsp("Captured HSP", captured_hsp);
      // Get reference pixel data from the memory and compute expected MSE
      expected_mse = new[hsid_x_top_gen.library_size];
      for (int j = 0; j < hsid_x_top_gen.library_size; j++) begin
        da_addr = hsid_x_top_gen.library_pixel_addr_w + (j * 4 * hsid_x_top_gen.hsp_bands_packs); // Address for each band
        expected_pixel_mem(da_addr, hsid_x_top_gen.hsp_bands, reference_hsp);
        hsid_x_top_gen.sq_df_acc_vctr(captured_hsp, reference_hsp, acc_int);
        hsid_x_top_gen.mse(acc_int, expected_mse[j], expected_mse_of[j]);
        hsid_x_top_gen.display_hsp("Reference HSP", reference_hsp);
        // $display("Accumulator: %p, MSE: %0d, Overflow: %0b", acc_int, expected_mse[j], expected_mse_of[j]);
        // $display("Library Pixel %0d: %p, MSE: %0d", j, reference_hsp, expected_mse[j]);
      end
      // $display(" - Vector sizes: captured %0d, reference %0d, accumulator %0d", captured_hsp.size(), reference_hsp.size(), acc_int.size());
      $display(" - Expected MSE values: %p", expected_mse);

      // Compute expected min and max MSE values and references
      hsid_x_top_gen.min_max_mse(expected_mse,
        min_mse_value_expected, max_mse_value_expected,
        min_mse_ref_expected, max_mse_ref_expected);

      $display(" - Expected min MSE: %0d, ref: %0d", min_mse_value_expected, min_mse_ref_expected);
      $display(" - Expected max MSE: %0d, ref: %0d", max_mse_value_expected, max_mse_ref_expected);

      // Initialize variables
      library_size_w = {{WORD_WIDTH-HSP_LIBRARY_WIDTH{1'b0}},hsid_x_top_gen.library_size};
      pixel_bands_w = {{WORD_WIDTH-HSP_BANDS_WIDTH{1'b0}}, hsid_x_top_gen.hsp_bands};
      captured_pixel_addr_w = hsid_x_top_gen.captured_pixel_addr_w;
      library_pixel_addr_w = hsid_x_top_gen.library_pixel_addr_w;

      // Check status register
      // assert_read_reg(HSID_X_CTRL_STATUS, STATUS_IDLE);

      // Initialize registers
      write_reg(reg_req, HSID_X_CTRL_CAPTURED_PIXEL_ADDR, captured_pixel_addr_w);
      write_reg(reg_req, HSID_X_CTRL_LIBRARY_PIXEL_ADDR, library_pixel_addr_w);
      write_reg(reg_req, HSID_X_CTRL_PIXEL_BANDS, pixel_bands_w);
      write_reg(reg_req, HSID_X_CTRL_LIBRARY_SIZE, library_size_w);


      // Check initialized values
      assert_read_reg(HSID_X_CTRL_LIBRARY_SIZE, library_size_w);
      assert_read_reg(HSID_X_CTRL_PIXEL_BANDS, pixel_bands_w);
      assert_read_reg(HSID_X_CTRL_CAPTURED_PIXEL_ADDR, captured_pixel_addr_w);
      assert_read_reg(HSID_X_CTRL_LIBRARY_PIXEL_ADDR, library_pixel_addr_w);

      // Start the processing
      write_reg(reg_req, HSID_X_CTRL_STATUS, STATUS_START);

      // Wait for the processing to complete, but add a delay to avoid problems with the clock
      wait (hsid_x_int_o == 1'b1);
      #8;
      assert_read_reg(HSID_X_CTRL_STATUS, STATUS_DONE);
      #10;
      assert_read_reg(HSID_X_CTRL_STATUS, STATUS_IDLE);

      // // Check the MSE results
      assert_read_reg(HSID_X_CTRL_MSE_MIN_REF, {{(WORD_WIDTH-HSP_LIBRARY_WIDTH){1'b0}}, min_mse_ref_expected });
      assert_read_reg(HSID_X_CTRL_MSE_MIN_VALUE, min_mse_value_expected);
      assert_read_reg(HSID_X_CTRL_MSE_MAX_REF, {{(WORD_WIDTH-HSP_LIBRARY_WIDTH){1'b0}}, max_mse_ref_expected });
      assert_read_reg(HSID_X_CTRL_MSE_MAX_VALUE, max_mse_value_expected);

      #20;

    end

    $finish;

  end

  always
    #5 clk = ! clk;

  // initial begin
  //   #20000; $finish; // Timeout if the test does not finish
  // end

  task assert_read_reg(input hsid_x_ctrl_id_e ctrl_id, logic [WORD_WIDTH-1:0] expected);
    read_reg(reg_req, ctrl_id);
    assert_value(reg_rsp.rdata, expected, $sformatf("BUS read addr: 0x%0h (%s)", addr_reg(ctrl_id), ctrl_id.name()));
  endtask

  task expected_pixel_mem(input logic [31:0] addr, input logic [HSP_BANDS_WIDTH-1:0] bands, output logic [DATA_WIDTH-1:0] hsp []);
    logic [DATA_WIDTH-1:0] msb_pixel_value;
    logic [DATA_WIDTH-1:0] lsb_pixel_value;
    hsp = new[bands];
    for (int i = 0; i < bands; i=i+2) begin
      msb_pixel_value = addr[WORD_WIDTH-1:DATA_WIDTH] & TEST_MEM_MASK;
      lsb_pixel_value = addr[DATA_WIDTH-1:0] & TEST_MEM_MASK;
      // $display("Reading pixel data from address: 0x%0h: 0x%0h", addr, masked_data);
      hsp[i] = lsb_pixel_value;
      hsp[i+1] = msb_pixel_value;
      addr = addr + 4;
    end
  endtask

endmodule